module s_box(
    input clk,
    input [7:0] inByte,
    output reg [7:0] subByte
);

// The whole s-box table
//reg [7:0] rijndael_sbox[255:0] = {8'h63, 8'h7C, 8'h77, 8'h7B, 8'hF2, 8'h6B, 8'h6F, 8'hC5, 8'h30, 8'h01, 8'h67, 8'h2B, 8'hFE, 8'hD7, 8'hAB, 8'h76, 8'hCA, 8'h82, 8'hC9, 8'h7D, 8'hFA, 8'h59, 8'h47, 8'hF0, 8'hAD, 8'hD4, 8'hA2, 8'hAF, 8'h9C, 8'hA4, 8'h72, 8'hC0, 8'hB7, 8'hFD, 8'h93, 8'h26, 8'h36, 8'h3F, 8'hF7, 8'hCC, 8'h34, 8'hA5, 8'hE5, 8'hF1, 8'h71, 8'hD8, 8'h31, 8'h15, 8'h04, 8'hC7, 8'h23, 8'hC3, 8'h18, 8'h96, 8'h05, 8'h9A, 8'h07, 8'h12, 8'h80, 8'hE2, 8'hEB, 8'h27, 8'hB2, 8'h75, 8'h09, 8'h83, 8'h2C, 8'h1A, 8'h1B, 8'h6E, 8'h5A, 8'hA0, 8'h52, 8'h3B, 8'hD6, 8'hB3, 8'h29, 8'hE3, 8'h2F, 8'h84, 8'h53, 8'hD1, 8'h00, 8'hED, 8'h20, 8'hFC, 8'hB1, 8'h5B, 8'h6A, 8'hCB, 8'hBE, 8'h39, 8'h4A, 8'h4C, 8'h58, 8'hCF, 8'hD0, 8'hEF, 8'hAA, 8'hFB, 8'h43, 8'h4D, 8'h33, 8'h85, 8'h45, 8'hF9, 8'h02, 8'h7F, 8'h50, 8'h3C, 8'h9F, 8'hA8, 8'h51, 8'hA3, 8'h40, 8'h8F, 8'h92, 8'h9D, 8'h38, 8'hF5, 8'hBC, 8'hB6, 8'hDA, 8'h21, 8'h10, 8'hFF, 8'hF3, 8'hD2, 8'hCD, 8'h0C, 8'h13, 8'hEC, 8'h5F, 8'h97, 8'h44, 8'h17, 8'hC4, 8'hA7, 8'h7E, 8'h3D, 8'h64, 8'h5D, 8'h19, 8'h73, 8'h60, 8'h81, 8'h4F, 8'hDC, 8'h22, 8'h2A, 8'h90, 8'h88, 8'h46, 8'hEE, 8'hB8, 8'h14, 8'hDE, 8'h5E, 8'h0B, 8'hDB, 8'hE0, 8'h32, 8'h3A, 8'h0A, 8'h49, 8'h06, 8'h24, 8'h5C, 8'hC2, 8'hD3, 8'hAC, 8'h62, 8'h91, 8'h95, 8'hE4, 8'h79, 8'hE7, 8'hC8, 8'h37, 8'h6D, 8'h8D, 8'hD5, 8'h4E, 8'hA9, 8'h6C, 8'h56, 8'hF4, 8'hEA, 8'h65, 8'h7A, 8'hAE, 8'h08, 8'hBA, 8'h78, 8'h25, 8'h2E, 8'h1C, 8'hA6, 8'hB4, 8'hC6, 8'hE8, 8'hDD, 8'h74, 8'h1F, 8'h4B, 8'hBD, 8'h8B, 8'h8A, 8'h70, 8'h3E, 8'hB5, 8'h66, 8'h48, 8'h03, 8'hF6, 8'h0E, 8'h61, 8'h35, 8'h57, 8'hB9, 8'h86, 8'hC1, 8'h1D, 8'h9E, 8'hE1, 8'hF8, 8'h98, 8'h11, 8'h69, 8'hD9, 8'h8E, 8'h94, 8'h9B, 8'h1E, 8'h87, 8'hE9, 8'hCE, 8'h55, 8'h28, 8'hDF, 8'h8C, 8'hA1, 8'h89, 8'h0D, 8'hBF, 8'hE6, 8'h42, 8'h68, 8'h41, 8'h99, 8'h2D, 8'h0F, 8'hB0, 8'h54, 8'hBB, 8'h16};

always @(posedge clk) begin
  case(inByte)
        8'd0: subByte = 8'h63;
        8'd1: subByte = 8'h7c;
        8'd2: subByte = 8'h77;
        8'd3: subByte = 8'h7b;
        8'd4: subByte = 8'hf2;
        8'd5: subByte = 8'h6b;
        8'd6: subByte = 8'h6f;
        8'd7: subByte = 8'hc5;
        8'd8: subByte = 8'h30;
        8'd9: subByte = 8'h01;
        8'd10: subByte = 8'h67;
        8'd11: subByte = 8'h2b;
        8'd12: subByte = 8'hfe;
        8'd13: subByte = 8'hd7;
        8'd14: subByte = 8'hab;
        8'd15: subByte = 8'h76;
        8'd16: subByte = 8'hca;
        8'd17: subByte = 8'h82;
        8'd18: subByte = 8'hc9;
        8'd19: subByte = 8'h7d;
        8'd20: subByte = 8'hfa;
        8'd21: subByte = 8'h59;
        8'd22: subByte = 8'h47;
        8'd23: subByte = 8'hf0;
        8'd24: subByte = 8'had;
        8'd25: subByte = 8'hd4;
        8'd26: subByte = 8'ha2;
        8'd27: subByte = 8'haf;
        8'd28: subByte = 8'h9c;
        8'd29: subByte = 8'ha4;
        8'd30: subByte = 8'h72;
        8'd31: subByte = 8'hc0;
        8'd32: subByte = 8'hb7;
        8'd33: subByte = 8'hfd;
        8'd34: subByte = 8'h93;
        8'd35: subByte = 8'h26;
        8'd36: subByte = 8'h36;
        8'd37: subByte = 8'h3f;
        8'd38: subByte = 8'hf7;
        8'd39: subByte = 8'hcc;
        8'd40: subByte = 8'h34;
        8'd41: subByte = 8'ha5;
        8'd42: subByte = 8'he5;
        8'd43: subByte = 8'hf1;
        8'd44: subByte = 8'h71;
        8'd45: subByte = 8'hd8;
        8'd46: subByte = 8'h31;
        8'd47: subByte = 8'h15;
        8'd48: subByte = 8'h04;
        8'd49: subByte = 8'hc7;
        8'd50: subByte = 8'h23;
        8'd51: subByte = 8'hc3;
        8'd52: subByte = 8'h18;
        8'd53: subByte = 8'h96;
        8'd54: subByte = 8'h05;
        8'd55: subByte = 8'h9a;
        8'd56: subByte = 8'h07;
        8'd57: subByte = 8'h12;
        8'd58: subByte = 8'h80;
        8'd59: subByte = 8'he2;
        8'd60: subByte = 8'heb;
        8'd61: subByte = 8'h27;
        8'd62: subByte = 8'hb2;
        8'd63: subByte = 8'h75;
        8'd64: subByte = 8'h09;
        8'd65: subByte = 8'h83;
        8'd66: subByte = 8'h2c;
        8'd67: subByte = 8'h1a;
        8'd68: subByte = 8'h1b;
        8'd69: subByte = 8'h6e;
        8'd70: subByte = 8'h5a;
        8'd71: subByte = 8'ha0;
        8'd72: subByte = 8'h52;
        8'd73: subByte = 8'h3b;
        8'd74: subByte = 8'hd6;
        8'd75: subByte = 8'hb3;
        8'd76: subByte = 8'h29;
        8'd77: subByte = 8'he3;
        8'd78: subByte = 8'h2f;
        8'd79: subByte = 8'h84;
        8'd80: subByte = 8'h53;
        8'd81: subByte = 8'hd1;
        8'd82: subByte = 8'h00;
        8'd83: subByte = 8'hed;
        8'd84: subByte = 8'h20;
        8'd85: subByte = 8'hfc;
        8'd86: subByte = 8'hb1;
        8'd87: subByte = 8'h5b;
        8'd88: subByte = 8'h6a;
        8'd89: subByte = 8'hcb;
        8'd90: subByte = 8'hbe;
        8'd91: subByte = 8'h39;
        8'd92: subByte = 8'h4a;
        8'd93: subByte = 8'h4c;
        8'd94: subByte = 8'h58;
        8'd95: subByte = 8'hcf;
        8'd96: subByte = 8'hd0;
        8'd97: subByte = 8'hef;
        8'd98: subByte = 8'haa;
        8'd99: subByte = 8'hfb;
        8'd100: subByte = 8'h43;
        8'd101: subByte = 8'h4d;
        8'd102: subByte = 8'h33;
        8'd103: subByte = 8'h85;
        8'd104: subByte = 8'h45;
        8'd105: subByte = 8'hf9;
        8'd106: subByte = 8'h02;
        8'd107: subByte = 8'h7f;
        8'd108: subByte = 8'h50;
        8'd109: subByte = 8'h3c;
        8'd110: subByte = 8'h9f;
        8'd111: subByte = 8'ha8;
        8'd112: subByte = 8'h51;
        8'd113: subByte = 8'ha3;
        8'd114: subByte = 8'h40;
        8'd115: subByte = 8'h8f;
        8'd116: subByte = 8'h92;
        8'd117: subByte = 8'h9d;
        8'd118: subByte = 8'h38;
        8'd119: subByte = 8'hf5;
        8'd120: subByte = 8'hbc;
        8'd121: subByte = 8'hb6;
        8'd122: subByte = 8'hda;
        8'd123: subByte = 8'h21;
        8'd124: subByte = 8'h10;
        8'd125: subByte = 8'hff;
        8'd126: subByte = 8'hf3;
        8'd127: subByte = 8'hd2;
        8'd128: subByte = 8'hcd;
        8'd129: subByte = 8'h0c;
        8'd130: subByte = 8'h13;
        8'd131: subByte = 8'hec;
        8'd132: subByte = 8'h5f;
        8'd133: subByte = 8'h97;
        8'd134: subByte = 8'h44;
        8'd135: subByte = 8'h17;
        8'd136: subByte = 8'hc4;
        8'd137: subByte = 8'ha7;
        8'd138: subByte = 8'h7e;
        8'd139: subByte = 8'h3d;
        8'd140: subByte = 8'h64;
        8'd141: subByte = 8'h5d;
        8'd142: subByte = 8'h19;
        8'd143: subByte = 8'h73;
        8'd144: subByte = 8'h60;
        8'd145: subByte = 8'h81;
        8'd146: subByte = 8'h4f;
        8'd147: subByte = 8'hdc;
        8'd148: subByte = 8'h22;
        8'd149: subByte = 8'h2a;
        8'd150: subByte = 8'h90;
        8'd151: subByte = 8'h88;
        8'd152: subByte = 8'h46;
        8'd153: subByte = 8'hee;
        8'd154: subByte = 8'hb8;
        8'd155: subByte = 8'h14;
        8'd156: subByte = 8'hde;
        8'd157: subByte = 8'h5e;
        8'd158: subByte = 8'h0b;
        8'd159: subByte = 8'hdb;
        8'd160: subByte = 8'he0;
        8'd161: subByte = 8'h32;
        8'd162: subByte = 8'h3a;
        8'd163: subByte = 8'h0a;
        8'd164: subByte = 8'h49;
        8'd165: subByte = 8'h06;
        8'd166: subByte = 8'h24;
        8'd167: subByte = 8'h5c;
        8'd168: subByte = 8'hc2;
        8'd169: subByte = 8'hd3;
        8'd170: subByte = 8'hac;
        8'd171: subByte = 8'h62;
        8'd172: subByte = 8'h91;
        8'd173: subByte = 8'h95;
        8'd174: subByte = 8'he4;
        8'd175: subByte = 8'h79;
        8'd176: subByte = 8'he7;
        8'd177: subByte = 8'hc8;
        8'd178: subByte = 8'h37;
        8'd179: subByte = 8'h6d;
        8'd180: subByte = 8'h8d;
        8'd181: subByte = 8'hd5;
        8'd182: subByte = 8'h4e;
        8'd183: subByte = 8'ha9;
        8'd184: subByte = 8'h6c;
        8'd185: subByte = 8'h56;
        8'd186: subByte = 8'hf4;
        8'd187: subByte = 8'hea;
        8'd188: subByte = 8'h65;
        8'd189: subByte = 8'h7a;
        8'd190: subByte = 8'hae;
        8'd191: subByte = 8'h08;
        8'd192: subByte = 8'hba;
        8'd193: subByte = 8'h78;
        8'd194: subByte = 8'h25;
        8'd195: subByte = 8'h2e;
        8'd196: subByte = 8'h1c;
        8'd197: subByte = 8'ha6;
        8'd198: subByte = 8'hb4;
        8'd199: subByte = 8'hc6;
        8'd200: subByte = 8'he8;
        8'd201: subByte = 8'hdd;
        8'd202: subByte = 8'h74;
        8'd203: subByte = 8'h1f;
        8'd204: subByte = 8'h4b;
        8'd205: subByte = 8'hbd;
        8'd206: subByte = 8'h8b;
        8'd207: subByte = 8'h8a;
        8'd208: subByte = 8'h70;
        8'd209: subByte = 8'h3e;
        8'd210: subByte = 8'hb5;
        8'd211: subByte = 8'h66;
        8'd212: subByte = 8'h48;
        8'd213: subByte = 8'h03;
        8'd214: subByte = 8'hf6;
        8'd215: subByte = 8'h0e;
        8'd216: subByte = 8'h61;
        8'd217: subByte = 8'h35;
        8'd218: subByte = 8'h57;
        8'd219: subByte = 8'hb9;
        8'd220: subByte = 8'h86;
        8'd221: subByte = 8'hc1;
        8'd222: subByte = 8'h1d;
        8'd223: subByte = 8'h9e;
        8'd224: subByte = 8'he1;
        8'd225: subByte = 8'hf8;
        8'd226: subByte = 8'h98;
        8'd227: subByte = 8'h11;
        8'd228: subByte = 8'h69;
        8'd229: subByte = 8'hd9;
        8'd230: subByte = 8'h8e;
        8'd231: subByte = 8'h94;
        8'd232: subByte = 8'h9b;
        8'd233: subByte = 8'h1e;
        8'd234: subByte = 8'h87;
        8'd235: subByte = 8'he9;
        8'd236: subByte = 8'hce;
        8'd237: subByte = 8'h55;
        8'd238: subByte = 8'h28;
        8'd239: subByte = 8'hdf;
        8'd240: subByte = 8'h8c;
        8'd241: subByte = 8'ha1;
        8'd242: subByte = 8'h89;
        8'd243: subByte = 8'h0d;
        8'd244: subByte = 8'hbf;
        8'd245: subByte = 8'he6;
        8'd246: subByte = 8'h42;
        8'd247: subByte = 8'h68;
        8'd248: subByte = 8'h41;
        8'd249: subByte = 8'h99;
        8'd250: subByte = 8'h2d;
        8'd251: subByte = 8'h0f;
        8'd252: subByte = 8'hb0;
        8'd253: subByte = 8'h54;
        8'd254: subByte = 8'hbb;
        8'd255: subByte = 8'h16;
  endcase
  //$display("index=%h, val=%h", inByte, subByte);
end

endmodule